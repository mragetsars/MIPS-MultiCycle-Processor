module Constant_1 (
    output [15:0] One
);
    assign One = 16'd1;
endmodule

module Constant_0 (
    output [15:0] Zero
);
    assign Zero = 16'd0;
endmodule