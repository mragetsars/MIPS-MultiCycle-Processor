module Adder16 (
    input  [15:0] A,
    input  [15:0] B,
    output [15:0] Sum
);
    assign Sum = A + B;
endmodule


